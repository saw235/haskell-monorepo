// Test file for minimal SystemVerilog parser
// This file contains valid SystemVerilog according to the minimal grammar

module simple_module;
endmodule

module counter;
endmodule

module memory_controller;
endmodule 